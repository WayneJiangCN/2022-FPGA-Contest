module CORES 
#( 
parameter CTRL_PORT_NUM     = 2,
parameter UJTAG_SEL         = 0,
parameter AREA_SPEED        = 0,    //0~5
parameter FLA0_MEM_STYLE         = 1,
parameter FLA0_TRIG_PORT_NUM     = 1,
parameter FLA0_MAX_SEQ_LEVEL     = 1,
parameter FLA0_EN_WINDOWS        = 0,
parameter FLA0_CLK_EDGE          = 1,
parameter FLA0_DATA_DEPTH        = 9,
parameter FLA0_EN_STOR_QUAL      = 0,
parameter FLA0_DATA_SAME_AS_TRIG = 1,
parameter FLA0_DATA_WIDTH        = 5,
parameter FLA0_TRIG0_PORT_WIDTH  = 5,
parameter FLA0_TRIG0_MATCH_UNIT  = 1,
parameter FLA0_TRIG0_CNT_WIDTH   = 0,
parameter FLA0_TRIG0_MATCH_TYPE  = 1,
parameter FLA0_TRIG0_EXCLUDE     = 0,
parameter FLA0_TRIG1_PORT_WIDTH  = 8,
parameter FLA0_TRIG1_MATCH_UNIT  = 1,
parameter FLA0_TRIG1_CNT_WIDTH   = 0,
parameter FLA0_TRIG1_MATCH_TYPE  = 1,
parameter FLA0_TRIG1_EXCLUDE     = 0,
parameter FLA0_TRIG2_PORT_WIDTH  = 8,
parameter FLA0_TRIG2_MATCH_UNIT  = 1,
parameter FLA0_TRIG2_CNT_WIDTH   = 0,
parameter FLA0_TRIG2_MATCH_TYPE  = 1,
parameter FLA0_TRIG2_EXCLUDE     = 0,
parameter FLA0_TRIG3_PORT_WIDTH  = 8,
parameter FLA0_TRIG3_MATCH_UNIT  = 1,
parameter FLA0_TRIG3_CNT_WIDTH   = 0,
parameter FLA0_TRIG3_MATCH_TYPE  = 1,
parameter FLA0_TRIG3_EXCLUDE     = 0,
parameter FLA0_TRIG4_PORT_WIDTH  = 8,
parameter FLA0_TRIG4_MATCH_UNIT  = 1,
parameter FLA0_TRIG4_CNT_WIDTH   = 0,
parameter FLA0_TRIG4_MATCH_TYPE  = 1,
parameter FLA0_TRIG4_EXCLUDE     = 0,
parameter FLA0_TRIG5_PORT_WIDTH  = 8,
parameter FLA0_TRIG5_MATCH_UNIT  = 1,
parameter FLA0_TRIG5_CNT_WIDTH   = 0,
parameter FLA0_TRIG5_MATCH_TYPE  = 1,
parameter FLA0_TRIG5_EXCLUDE     = 0,
parameter FLA0_TRIG6_PORT_WIDTH  = 8,
parameter FLA0_TRIG6_MATCH_UNIT  = 1,
parameter FLA0_TRIG6_CNT_WIDTH   = 0,
parameter FLA0_TRIG6_MATCH_TYPE  = 1,
parameter FLA0_TRIG6_EXCLUDE     = 0,
parameter FLA0_TRIG7_PORT_WIDTH  = 8,
parameter FLA0_TRIG7_MATCH_UNIT  = 1,
parameter FLA0_TRIG7_CNT_WIDTH   = 0,
parameter FLA0_TRIG7_MATCH_TYPE  = 1,
parameter FLA0_TRIG7_EXCLUDE     = 0,
parameter FLA0_TRIG8_PORT_WIDTH  = 8,
parameter FLA0_TRIG8_MATCH_UNIT  = 1,
parameter FLA0_TRIG8_CNT_WIDTH   = 0,
parameter FLA0_TRIG8_MATCH_TYPE  = 1,
parameter FLA0_TRIG8_EXCLUDE     = 0,
parameter FLA0_TRIG9_PORT_WIDTH  = 8,
parameter FLA0_TRIG9_MATCH_UNIT  = 1,
parameter FLA0_TRIG9_CNT_WIDTH   = 0,
parameter FLA0_TRIG9_MATCH_TYPE  = 1,
parameter FLA0_TRIG9_EXCLUDE     = 0,
parameter FLA0_TRIG10_PORT_WIDTH  = 8,
parameter FLA0_TRIG10_MATCH_UNIT  = 1,
parameter FLA0_TRIG10_CNT_WIDTH   = 0,
parameter FLA0_TRIG10_MATCH_TYPE  = 1,
parameter FLA0_TRIG10_EXCLUDE     = 0,
parameter FLA0_TRIG11_PORT_WIDTH  = 8,
parameter FLA0_TRIG11_MATCH_UNIT  = 1,
parameter FLA0_TRIG11_CNT_WIDTH   = 0,
parameter FLA0_TRIG11_MATCH_TYPE  = 1,
parameter FLA0_TRIG11_EXCLUDE     = 0,
parameter FLA0_TRIG12_PORT_WIDTH  = 8,
parameter FLA0_TRIG12_MATCH_UNIT  = 1,
parameter FLA0_TRIG12_CNT_WIDTH   = 0,
parameter FLA0_TRIG12_MATCH_TYPE  = 1,
parameter FLA0_TRIG12_EXCLUDE     = 0,
parameter FLA0_TRIG13_PORT_WIDTH  = 8,
parameter FLA0_TRIG13_MATCH_UNIT  = 1,
parameter FLA0_TRIG13_CNT_WIDTH   = 0,
parameter FLA0_TRIG13_MATCH_TYPE  = 1,
parameter FLA0_TRIG13_EXCLUDE     = 0,
parameter FLA0_TRIG14_PORT_WIDTH  = 8,
parameter FLA0_TRIG14_MATCH_UNIT  = 1,
parameter FLA0_TRIG14_CNT_WIDTH   = 0,
parameter FLA0_TRIG14_MATCH_TYPE  = 1,
parameter FLA0_TRIG14_EXCLUDE     = 0,
parameter FLA0_TRIG15_PORT_WIDTH  = 8,
parameter FLA0_TRIG15_MATCH_UNIT  = 1,
parameter FLA0_TRIG15_CNT_WIDTH   = 0,
parameter FLA0_TRIG15_MATCH_TYPE  = 1,
parameter FLA0_TRIG15_EXCLUDE     = 0,
parameter FLA1_MEM_STYLE         = 1,
parameter FLA1_TRIG_PORT_NUM     = 1,
parameter FLA1_MAX_SEQ_LEVEL     = 1,
parameter FLA1_EN_WINDOWS        = 0,
parameter FLA1_CLK_EDGE          = 1,
parameter FLA1_DATA_DEPTH        = 9,
parameter FLA1_EN_STOR_QUAL      = 0,
parameter FLA1_DATA_SAME_AS_TRIG = 1,
parameter FLA1_DATA_WIDTH        = 24,
parameter FLA1_TRIG0_PORT_WIDTH  = 24,
parameter FLA1_TRIG0_MATCH_UNIT  = 1,
parameter FLA1_TRIG0_CNT_WIDTH   = 0,
parameter FLA1_TRIG0_MATCH_TYPE  = 1,
parameter FLA1_TRIG0_EXCLUDE     = 0,
parameter FLA1_TRIG1_PORT_WIDTH  = 8,
parameter FLA1_TRIG1_MATCH_UNIT  = 1,
parameter FLA1_TRIG1_CNT_WIDTH   = 0,
parameter FLA1_TRIG1_MATCH_TYPE  = 1,
parameter FLA1_TRIG1_EXCLUDE     = 0,
parameter FLA1_TRIG2_PORT_WIDTH  = 8,
parameter FLA1_TRIG2_MATCH_UNIT  = 1,
parameter FLA1_TRIG2_CNT_WIDTH   = 0,
parameter FLA1_TRIG2_MATCH_TYPE  = 1,
parameter FLA1_TRIG2_EXCLUDE     = 0,
parameter FLA1_TRIG3_PORT_WIDTH  = 8,
parameter FLA1_TRIG3_MATCH_UNIT  = 1,
parameter FLA1_TRIG3_CNT_WIDTH   = 0,
parameter FLA1_TRIG3_MATCH_TYPE  = 1,
parameter FLA1_TRIG3_EXCLUDE     = 0,
parameter FLA1_TRIG4_PORT_WIDTH  = 8,
parameter FLA1_TRIG4_MATCH_UNIT  = 1,
parameter FLA1_TRIG4_CNT_WIDTH   = 0,
parameter FLA1_TRIG4_MATCH_TYPE  = 1,
parameter FLA1_TRIG4_EXCLUDE     = 0,
parameter FLA1_TRIG5_PORT_WIDTH  = 8,
parameter FLA1_TRIG5_MATCH_UNIT  = 1,
parameter FLA1_TRIG5_CNT_WIDTH   = 0,
parameter FLA1_TRIG5_MATCH_TYPE  = 1,
parameter FLA1_TRIG5_EXCLUDE     = 0,
parameter FLA1_TRIG6_PORT_WIDTH  = 8,
parameter FLA1_TRIG6_MATCH_UNIT  = 1,
parameter FLA1_TRIG6_CNT_WIDTH   = 0,
parameter FLA1_TRIG6_MATCH_TYPE  = 1,
parameter FLA1_TRIG6_EXCLUDE     = 0,
parameter FLA1_TRIG7_PORT_WIDTH  = 8,
parameter FLA1_TRIG7_MATCH_UNIT  = 1,
parameter FLA1_TRIG7_CNT_WIDTH   = 0,
parameter FLA1_TRIG7_MATCH_TYPE  = 1,
parameter FLA1_TRIG7_EXCLUDE     = 0,
parameter FLA1_TRIG8_PORT_WIDTH  = 8,
parameter FLA1_TRIG8_MATCH_UNIT  = 1,
parameter FLA1_TRIG8_CNT_WIDTH   = 0,
parameter FLA1_TRIG8_MATCH_TYPE  = 1,
parameter FLA1_TRIG8_EXCLUDE     = 0,
parameter FLA1_TRIG9_PORT_WIDTH  = 8,
parameter FLA1_TRIG9_MATCH_UNIT  = 1,
parameter FLA1_TRIG9_CNT_WIDTH   = 0,
parameter FLA1_TRIG9_MATCH_TYPE  = 1,
parameter FLA1_TRIG9_EXCLUDE     = 0,
parameter FLA1_TRIG10_PORT_WIDTH  = 8,
parameter FLA1_TRIG10_MATCH_UNIT  = 1,
parameter FLA1_TRIG10_CNT_WIDTH   = 0,
parameter FLA1_TRIG10_MATCH_TYPE  = 1,
parameter FLA1_TRIG10_EXCLUDE     = 0,
parameter FLA1_TRIG11_PORT_WIDTH  = 8,
parameter FLA1_TRIG11_MATCH_UNIT  = 1,
parameter FLA1_TRIG11_CNT_WIDTH   = 0,
parameter FLA1_TRIG11_MATCH_TYPE  = 1,
parameter FLA1_TRIG11_EXCLUDE     = 0,
parameter FLA1_TRIG12_PORT_WIDTH  = 8,
parameter FLA1_TRIG12_MATCH_UNIT  = 1,
parameter FLA1_TRIG12_CNT_WIDTH   = 0,
parameter FLA1_TRIG12_MATCH_TYPE  = 1,
parameter FLA1_TRIG12_EXCLUDE     = 0,
parameter FLA1_TRIG13_PORT_WIDTH  = 8,
parameter FLA1_TRIG13_MATCH_UNIT  = 1,
parameter FLA1_TRIG13_CNT_WIDTH   = 0,
parameter FLA1_TRIG13_MATCH_TYPE  = 1,
parameter FLA1_TRIG13_EXCLUDE     = 0,
parameter FLA1_TRIG14_PORT_WIDTH  = 8,
parameter FLA1_TRIG14_MATCH_UNIT  = 1,
parameter FLA1_TRIG14_CNT_WIDTH   = 0,
parameter FLA1_TRIG14_MATCH_TYPE  = 1,
parameter FLA1_TRIG14_EXCLUDE     = 0,
parameter FLA1_TRIG15_PORT_WIDTH  = 8,
parameter FLA1_TRIG15_MATCH_UNIT  = 1,
parameter FLA1_TRIG15_CNT_WIDTH   = 0,
parameter FLA1_TRIG15_MATCH_TYPE  = 1,
parameter FLA1_TRIG15_EXCLUDE     = 0
) ( 
input  dbc_urck_in,                 //TCK from user pad 
input  dbc_utdi_in,                 //TDI from user pad 
input  [FLA0_DATA_WIDTH-1:0]  fla0_data_i, 
input  [FLA0_TRIG0_PORT_WIDTH-1:0] fla0_trig0_i, 
input  [FLA0_TRIG1_PORT_WIDTH-1:0] fla0_trig1_i, 
input  [FLA0_TRIG2_PORT_WIDTH-1:0] fla0_trig2_i, 
input  [FLA0_TRIG3_PORT_WIDTH-1:0] fla0_trig3_i, 
input  [FLA0_TRIG4_PORT_WIDTH-1:0] fla0_trig4_i, 
input  [FLA0_TRIG5_PORT_WIDTH-1:0] fla0_trig5_i, 
input  [FLA0_TRIG6_PORT_WIDTH-1:0] fla0_trig6_i, 
input  [FLA0_TRIG7_PORT_WIDTH-1:0] fla0_trig7_i, 
input  [FLA0_TRIG8_PORT_WIDTH-1:0] fla0_trig8_i, 
input  [FLA0_TRIG9_PORT_WIDTH-1:0] fla0_trig9_i, 
input  [FLA0_TRIG10_PORT_WIDTH-1:0] fla0_trig10_i, 
input  [FLA0_TRIG11_PORT_WIDTH-1:0] fla0_trig11_i, 
input  [FLA0_TRIG12_PORT_WIDTH-1:0] fla0_trig12_i, 
input  [FLA0_TRIG13_PORT_WIDTH-1:0] fla0_trig13_i, 
input  [FLA0_TRIG14_PORT_WIDTH-1:0] fla0_trig14_i, 
input  [FLA0_TRIG15_PORT_WIDTH-1:0] fla0_trig15_i, 
input fla0_rstn , 
input fla0_clk , 
input  [FLA1_DATA_WIDTH-1:0]  fla1_data_i, 
input  [FLA1_TRIG0_PORT_WIDTH-1:0] fla1_trig0_i, 
input  [FLA1_TRIG1_PORT_WIDTH-1:0] fla1_trig1_i, 
input  [FLA1_TRIG2_PORT_WIDTH-1:0] fla1_trig2_i, 
input  [FLA1_TRIG3_PORT_WIDTH-1:0] fla1_trig3_i, 
input  [FLA1_TRIG4_PORT_WIDTH-1:0] fla1_trig4_i, 
input  [FLA1_TRIG5_PORT_WIDTH-1:0] fla1_trig5_i, 
input  [FLA1_TRIG6_PORT_WIDTH-1:0] fla1_trig6_i, 
input  [FLA1_TRIG7_PORT_WIDTH-1:0] fla1_trig7_i, 
input  [FLA1_TRIG8_PORT_WIDTH-1:0] fla1_trig8_i, 
input  [FLA1_TRIG9_PORT_WIDTH-1:0] fla1_trig9_i, 
input  [FLA1_TRIG10_PORT_WIDTH-1:0] fla1_trig10_i, 
input  [FLA1_TRIG11_PORT_WIDTH-1:0] fla1_trig11_i, 
input  [FLA1_TRIG12_PORT_WIDTH-1:0] fla1_trig12_i, 
input  [FLA1_TRIG13_PORT_WIDTH-1:0] fla1_trig13_i, 
input  [FLA1_TRIG14_PORT_WIDTH-1:0] fla1_trig14_i, 
input  [FLA1_TRIG15_PORT_WIDTH-1:0] fla1_trig15_i, 
input fla1_rstn , 
input fla1_clk
)/* synthesis syn_noprune = 1 */;
wire capture_wire,drck1_wire, reset_wire,sel1_wire,shift_wire,update_wire,tdi_wire,tdo1_wire;
GTP_SCANCHAIN_E1 #( 
.CHAIN_NUM  (1)
)
 u_GTP_SCANCHAIN_PG (
                    .CAPDR(capture_wire),
                    .TCK_USER(drck1_wire),
                    .RST(reset_wire),
                    .FLG_USER(sel1_wire),
                    .SHFTDR(shift_wire),
                    .TDI_USER(tdi_wire),
                    .UPDR(update_wire),
                    .TDO_USER(tdo1_wire)
                    )/* synthesis syn_noprune = 1*/;
 wire drck_o;  
wire conf_tdi;  
wire [15:0] conf_sel;  
wire [4:0] id_o;  
wire [15:0] hub_tdo;  
wire capt_o;  
wire shift_d;
ips_jtag_hub_v1_3 
#( 
.CTRL_PORT_NUM  (CTRL_PORT_NUM),         //the number of usr_app connect with jtag_hub
.UJTAG_SEL      (UJTAG_SEL)              //1:use jtagif ;0:use scanchain
)
u_jtag_hub(
// for USER JTAGIF
.urck_in       (dbc_urck_in),                  //TCK from user pad 
.utdi_in       (dbc_utdi_in),                  //TDI from user pad 
// for JTAG_interface    
.tdi_in       (tdi_wire),                 //TDI for user data register;
.tdo_out      (tdo1_wire),                //TDO for user data register 
.reset_dr     (reset_wire),               //active high reset when TAP state in e_TEST_LOGIC_RESET state
.shift_in     (shift_wire),              //TAP state in e_SHIFT_DR,for pg30 design is reversed
.update_in    (update_wire),              //TAP state in e_UPDATE_DR
.capture_in   (capture_wire),             //TAP state in e_CAPTURE_DR
.sel_in       (sel1_wire),                 //user data register is selected
.h_rstn       (1'b1),.drck_in      (drck1_wire),                //TCK for user data register
// for user_app interface(debug_core,etc)
.drck_o       (drck_o),                //transfer TCK to each user_app
.conf_tdi     (conf_tdi),              //transfer TDI to each user_app
.conf_sel     (conf_sel),              //select config module which indicated by ID
.id_o         (id_o),                  //ID number indication
.capt_o       (capt_o),                 //capture
.hub_tdo      (hub_tdo),                //read back signal from each user_app
.shift_d      (shift_d)
)/* synthesis syn_noprune = 1*/; 
ips_dbc_debug_core_v1_4 
#( 
.AREA_SPEED           (AREA_SPEED), 
.MEM_STYLE            (FLA0_MEM_STYLE), 
.TRIG_PORT_NUM        (FLA0_TRIG_PORT_NUM), 
.MAX_SEQ_LEVEL        (FLA0_MAX_SEQ_LEVEL), 
.EN_WINDOWS           (FLA0_EN_WINDOWS),
.CLK_EDGE             (FLA0_CLK_EDGE), 
.DATA_DEPTH           (FLA0_DATA_DEPTH), 
.EN_STOR_QUAL         (FLA0_EN_STOR_QUAL), 
.DATA_SAME_AS_TRIG    (FLA0_DATA_SAME_AS_TRIG), 
.DATA_WIDTH           (FLA0_DATA_WIDTH), 
.TRIG0_PORT_WIDTH           (FLA0_TRIG0_PORT_WIDTH ), 
.TRIG0_MATCH_UNIT            (FLA0_TRIG0_MATCH_UNIT ), 
.TRIG0_CNT_WIDTH           (FLA0_TRIG0_CNT_WIDTH ), 
.TRIG0_MATCH_TYPE           (FLA0_TRIG0_MATCH_TYPE ), 
.TRIG0_EXCLUDE           (FLA0_TRIG0_EXCLUDE ), 
.TRIG1_PORT_WIDTH           (FLA0_TRIG1_PORT_WIDTH ), 
.TRIG1_MATCH_UNIT            (FLA0_TRIG1_MATCH_UNIT ), 
.TRIG1_CNT_WIDTH           (FLA0_TRIG1_CNT_WIDTH ), 
.TRIG1_MATCH_TYPE           (FLA0_TRIG1_MATCH_TYPE ), 
.TRIG1_EXCLUDE           (FLA0_TRIG1_EXCLUDE ), 
.TRIG2_PORT_WIDTH           (FLA0_TRIG2_PORT_WIDTH ), 
.TRIG2_MATCH_UNIT            (FLA0_TRIG2_MATCH_UNIT ), 
.TRIG2_CNT_WIDTH           (FLA0_TRIG2_CNT_WIDTH ), 
.TRIG2_MATCH_TYPE           (FLA0_TRIG2_MATCH_TYPE ), 
.TRIG2_EXCLUDE           (FLA0_TRIG2_EXCLUDE ), 
.TRIG3_PORT_WIDTH           (FLA0_TRIG3_PORT_WIDTH ), 
.TRIG3_MATCH_UNIT            (FLA0_TRIG3_MATCH_UNIT ), 
.TRIG3_CNT_WIDTH           (FLA0_TRIG3_CNT_WIDTH ), 
.TRIG3_MATCH_TYPE           (FLA0_TRIG3_MATCH_TYPE ), 
.TRIG3_EXCLUDE           (FLA0_TRIG3_EXCLUDE ), 
.TRIG4_PORT_WIDTH           (FLA0_TRIG4_PORT_WIDTH ), 
.TRIG4_MATCH_UNIT            (FLA0_TRIG4_MATCH_UNIT ), 
.TRIG4_CNT_WIDTH           (FLA0_TRIG4_CNT_WIDTH ), 
.TRIG4_MATCH_TYPE           (FLA0_TRIG4_MATCH_TYPE ), 
.TRIG4_EXCLUDE           (FLA0_TRIG4_EXCLUDE ), 
.TRIG5_PORT_WIDTH           (FLA0_TRIG5_PORT_WIDTH ), 
.TRIG5_MATCH_UNIT            (FLA0_TRIG5_MATCH_UNIT ), 
.TRIG5_CNT_WIDTH           (FLA0_TRIG5_CNT_WIDTH ), 
.TRIG5_MATCH_TYPE           (FLA0_TRIG5_MATCH_TYPE ), 
.TRIG5_EXCLUDE           (FLA0_TRIG5_EXCLUDE ), 
.TRIG6_PORT_WIDTH           (FLA0_TRIG6_PORT_WIDTH ), 
.TRIG6_MATCH_UNIT            (FLA0_TRIG6_MATCH_UNIT ), 
.TRIG6_CNT_WIDTH           (FLA0_TRIG6_CNT_WIDTH ), 
.TRIG6_MATCH_TYPE           (FLA0_TRIG6_MATCH_TYPE ), 
.TRIG6_EXCLUDE           (FLA0_TRIG6_EXCLUDE ), 
.TRIG7_PORT_WIDTH           (FLA0_TRIG7_PORT_WIDTH ), 
.TRIG7_MATCH_UNIT            (FLA0_TRIG7_MATCH_UNIT ), 
.TRIG7_CNT_WIDTH           (FLA0_TRIG7_CNT_WIDTH ), 
.TRIG7_MATCH_TYPE           (FLA0_TRIG7_MATCH_TYPE ), 
.TRIG7_EXCLUDE           (FLA0_TRIG7_EXCLUDE ), 
.TRIG8_PORT_WIDTH           (FLA0_TRIG8_PORT_WIDTH ), 
.TRIG8_MATCH_UNIT            (FLA0_TRIG8_MATCH_UNIT ), 
.TRIG8_CNT_WIDTH           (FLA0_TRIG8_CNT_WIDTH ), 
.TRIG8_MATCH_TYPE           (FLA0_TRIG8_MATCH_TYPE ), 
.TRIG8_EXCLUDE           (FLA0_TRIG8_EXCLUDE ), 
.TRIG9_PORT_WIDTH           (FLA0_TRIG9_PORT_WIDTH ), 
.TRIG9_MATCH_UNIT            (FLA0_TRIG9_MATCH_UNIT ), 
.TRIG9_CNT_WIDTH           (FLA0_TRIG9_CNT_WIDTH ), 
.TRIG9_MATCH_TYPE           (FLA0_TRIG9_MATCH_TYPE ), 
.TRIG9_EXCLUDE           (FLA0_TRIG9_EXCLUDE ), 
.TRIG10_PORT_WIDTH           (FLA0_TRIG10_PORT_WIDTH ), 
.TRIG10_MATCH_UNIT            (FLA0_TRIG10_MATCH_UNIT ), 
.TRIG10_CNT_WIDTH           (FLA0_TRIG10_CNT_WIDTH ), 
.TRIG10_MATCH_TYPE           (FLA0_TRIG10_MATCH_TYPE ), 
.TRIG10_EXCLUDE           (FLA0_TRIG10_EXCLUDE ), 
.TRIG11_PORT_WIDTH           (FLA0_TRIG11_PORT_WIDTH ), 
.TRIG11_MATCH_UNIT            (FLA0_TRIG11_MATCH_UNIT ), 
.TRIG11_CNT_WIDTH           (FLA0_TRIG11_CNT_WIDTH ), 
.TRIG11_MATCH_TYPE           (FLA0_TRIG11_MATCH_TYPE ), 
.TRIG11_EXCLUDE           (FLA0_TRIG11_EXCLUDE ), 
.TRIG12_PORT_WIDTH           (FLA0_TRIG12_PORT_WIDTH ), 
.TRIG12_MATCH_UNIT            (FLA0_TRIG12_MATCH_UNIT ), 
.TRIG12_CNT_WIDTH           (FLA0_TRIG12_CNT_WIDTH ), 
.TRIG12_MATCH_TYPE           (FLA0_TRIG12_MATCH_TYPE ), 
.TRIG12_EXCLUDE           (FLA0_TRIG12_EXCLUDE ), 
.TRIG13_PORT_WIDTH           (FLA0_TRIG13_PORT_WIDTH ), 
.TRIG13_MATCH_UNIT            (FLA0_TRIG13_MATCH_UNIT ), 
.TRIG13_CNT_WIDTH           (FLA0_TRIG13_CNT_WIDTH ), 
.TRIG13_MATCH_TYPE           (FLA0_TRIG13_MATCH_TYPE ), 
.TRIG13_EXCLUDE           (FLA0_TRIG13_EXCLUDE ), 
.TRIG14_PORT_WIDTH           (FLA0_TRIG14_PORT_WIDTH ), 
.TRIG14_MATCH_UNIT            (FLA0_TRIG14_MATCH_UNIT ), 
.TRIG14_CNT_WIDTH           (FLA0_TRIG14_CNT_WIDTH ), 
.TRIG14_MATCH_TYPE           (FLA0_TRIG14_MATCH_TYPE ), 
.TRIG14_EXCLUDE           (FLA0_TRIG14_EXCLUDE ), 
.TRIG15_PORT_WIDTH           (FLA0_TRIG15_PORT_WIDTH ), 
.TRIG15_MATCH_UNIT            (FLA0_TRIG15_MATCH_UNIT ), 
.TRIG15_CNT_WIDTH           (FLA0_TRIG15_CNT_WIDTH ), 
.TRIG15_MATCH_TYPE           (FLA0_TRIG15_MATCH_TYPE ), 
.TRIG15_EXCLUDE           (FLA0_TRIG15_EXCLUDE )
) 
u_debug_core_0( 
.drck_in      (drck_o),  
.hub_tdi      (conf_tdi),  
.id_i         (id_o),  
.shift_i      (shift_d), 
.capt_i               (capt_o),  
.conf_sel     (conf_sel[0]),  
.hub_tdo      (hub_tdo[0]),  
.clk          (fla0_clk),  
.resetn_i     (fla0_rstn),  
.trig0_i       (fla0_trig0_i),  
.trig1_i       (fla0_trig1_i),  
.trig2_i       (fla0_trig2_i),  
.trig3_i       (fla0_trig3_i),  
.trig4_i       (fla0_trig4_i),  
.trig5_i       (fla0_trig5_i),  
.trig6_i       (fla0_trig6_i),  
.trig7_i       (fla0_trig7_i),  
.trig8_i       (fla0_trig8_i),  
.trig9_i       (fla0_trig9_i),  
.trig10_i       (fla0_trig10_i),  
.trig11_i       (fla0_trig11_i),  
.trig12_i       (fla0_trig12_i),  
.trig13_i       (fla0_trig13_i),  
.trig14_i       (fla0_trig14_i),  
.trig15_i       (fla0_trig15_i),  
.data_i       (fla0_data_i)  
); 
ips_dbc_debug_core_v1_4 
#( 
.AREA_SPEED           (AREA_SPEED), 
.MEM_STYLE            (FLA1_MEM_STYLE), 
.TRIG_PORT_NUM        (FLA1_TRIG_PORT_NUM), 
.MAX_SEQ_LEVEL        (FLA1_MAX_SEQ_LEVEL), 
.EN_WINDOWS           (FLA1_EN_WINDOWS),
.CLK_EDGE             (FLA1_CLK_EDGE), 
.DATA_DEPTH           (FLA1_DATA_DEPTH), 
.EN_STOR_QUAL         (FLA1_EN_STOR_QUAL), 
.DATA_SAME_AS_TRIG    (FLA1_DATA_SAME_AS_TRIG), 
.DATA_WIDTH           (FLA1_DATA_WIDTH), 
.TRIG0_PORT_WIDTH           (FLA1_TRIG0_PORT_WIDTH ), 
.TRIG0_MATCH_UNIT            (FLA1_TRIG0_MATCH_UNIT ), 
.TRIG0_CNT_WIDTH           (FLA1_TRIG0_CNT_WIDTH ), 
.TRIG0_MATCH_TYPE           (FLA1_TRIG0_MATCH_TYPE ), 
.TRIG0_EXCLUDE           (FLA1_TRIG0_EXCLUDE ), 
.TRIG1_PORT_WIDTH           (FLA1_TRIG1_PORT_WIDTH ), 
.TRIG1_MATCH_UNIT            (FLA1_TRIG1_MATCH_UNIT ), 
.TRIG1_CNT_WIDTH           (FLA1_TRIG1_CNT_WIDTH ), 
.TRIG1_MATCH_TYPE           (FLA1_TRIG1_MATCH_TYPE ), 
.TRIG1_EXCLUDE           (FLA1_TRIG1_EXCLUDE ), 
.TRIG2_PORT_WIDTH           (FLA1_TRIG2_PORT_WIDTH ), 
.TRIG2_MATCH_UNIT            (FLA1_TRIG2_MATCH_UNIT ), 
.TRIG2_CNT_WIDTH           (FLA1_TRIG2_CNT_WIDTH ), 
.TRIG2_MATCH_TYPE           (FLA1_TRIG2_MATCH_TYPE ), 
.TRIG2_EXCLUDE           (FLA1_TRIG2_EXCLUDE ), 
.TRIG3_PORT_WIDTH           (FLA1_TRIG3_PORT_WIDTH ), 
.TRIG3_MATCH_UNIT            (FLA1_TRIG3_MATCH_UNIT ), 
.TRIG3_CNT_WIDTH           (FLA1_TRIG3_CNT_WIDTH ), 
.TRIG3_MATCH_TYPE           (FLA1_TRIG3_MATCH_TYPE ), 
.TRIG3_EXCLUDE           (FLA1_TRIG3_EXCLUDE ), 
.TRIG4_PORT_WIDTH           (FLA1_TRIG4_PORT_WIDTH ), 
.TRIG4_MATCH_UNIT            (FLA1_TRIG4_MATCH_UNIT ), 
.TRIG4_CNT_WIDTH           (FLA1_TRIG4_CNT_WIDTH ), 
.TRIG4_MATCH_TYPE           (FLA1_TRIG4_MATCH_TYPE ), 
.TRIG4_EXCLUDE           (FLA1_TRIG4_EXCLUDE ), 
.TRIG5_PORT_WIDTH           (FLA1_TRIG5_PORT_WIDTH ), 
.TRIG5_MATCH_UNIT            (FLA1_TRIG5_MATCH_UNIT ), 
.TRIG5_CNT_WIDTH           (FLA1_TRIG5_CNT_WIDTH ), 
.TRIG5_MATCH_TYPE           (FLA1_TRIG5_MATCH_TYPE ), 
.TRIG5_EXCLUDE           (FLA1_TRIG5_EXCLUDE ), 
.TRIG6_PORT_WIDTH           (FLA1_TRIG6_PORT_WIDTH ), 
.TRIG6_MATCH_UNIT            (FLA1_TRIG6_MATCH_UNIT ), 
.TRIG6_CNT_WIDTH           (FLA1_TRIG6_CNT_WIDTH ), 
.TRIG6_MATCH_TYPE           (FLA1_TRIG6_MATCH_TYPE ), 
.TRIG6_EXCLUDE           (FLA1_TRIG6_EXCLUDE ), 
.TRIG7_PORT_WIDTH           (FLA1_TRIG7_PORT_WIDTH ), 
.TRIG7_MATCH_UNIT            (FLA1_TRIG7_MATCH_UNIT ), 
.TRIG7_CNT_WIDTH           (FLA1_TRIG7_CNT_WIDTH ), 
.TRIG7_MATCH_TYPE           (FLA1_TRIG7_MATCH_TYPE ), 
.TRIG7_EXCLUDE           (FLA1_TRIG7_EXCLUDE ), 
.TRIG8_PORT_WIDTH           (FLA1_TRIG8_PORT_WIDTH ), 
.TRIG8_MATCH_UNIT            (FLA1_TRIG8_MATCH_UNIT ), 
.TRIG8_CNT_WIDTH           (FLA1_TRIG8_CNT_WIDTH ), 
.TRIG8_MATCH_TYPE           (FLA1_TRIG8_MATCH_TYPE ), 
.TRIG8_EXCLUDE           (FLA1_TRIG8_EXCLUDE ), 
.TRIG9_PORT_WIDTH           (FLA1_TRIG9_PORT_WIDTH ), 
.TRIG9_MATCH_UNIT            (FLA1_TRIG9_MATCH_UNIT ), 
.TRIG9_CNT_WIDTH           (FLA1_TRIG9_CNT_WIDTH ), 
.TRIG9_MATCH_TYPE           (FLA1_TRIG9_MATCH_TYPE ), 
.TRIG9_EXCLUDE           (FLA1_TRIG9_EXCLUDE ), 
.TRIG10_PORT_WIDTH           (FLA1_TRIG10_PORT_WIDTH ), 
.TRIG10_MATCH_UNIT            (FLA1_TRIG10_MATCH_UNIT ), 
.TRIG10_CNT_WIDTH           (FLA1_TRIG10_CNT_WIDTH ), 
.TRIG10_MATCH_TYPE           (FLA1_TRIG10_MATCH_TYPE ), 
.TRIG10_EXCLUDE           (FLA1_TRIG10_EXCLUDE ), 
.TRIG11_PORT_WIDTH           (FLA1_TRIG11_PORT_WIDTH ), 
.TRIG11_MATCH_UNIT            (FLA1_TRIG11_MATCH_UNIT ), 
.TRIG11_CNT_WIDTH           (FLA1_TRIG11_CNT_WIDTH ), 
.TRIG11_MATCH_TYPE           (FLA1_TRIG11_MATCH_TYPE ), 
.TRIG11_EXCLUDE           (FLA1_TRIG11_EXCLUDE ), 
.TRIG12_PORT_WIDTH           (FLA1_TRIG12_PORT_WIDTH ), 
.TRIG12_MATCH_UNIT            (FLA1_TRIG12_MATCH_UNIT ), 
.TRIG12_CNT_WIDTH           (FLA1_TRIG12_CNT_WIDTH ), 
.TRIG12_MATCH_TYPE           (FLA1_TRIG12_MATCH_TYPE ), 
.TRIG12_EXCLUDE           (FLA1_TRIG12_EXCLUDE ), 
.TRIG13_PORT_WIDTH           (FLA1_TRIG13_PORT_WIDTH ), 
.TRIG13_MATCH_UNIT            (FLA1_TRIG13_MATCH_UNIT ), 
.TRIG13_CNT_WIDTH           (FLA1_TRIG13_CNT_WIDTH ), 
.TRIG13_MATCH_TYPE           (FLA1_TRIG13_MATCH_TYPE ), 
.TRIG13_EXCLUDE           (FLA1_TRIG13_EXCLUDE ), 
.TRIG14_PORT_WIDTH           (FLA1_TRIG14_PORT_WIDTH ), 
.TRIG14_MATCH_UNIT            (FLA1_TRIG14_MATCH_UNIT ), 
.TRIG14_CNT_WIDTH           (FLA1_TRIG14_CNT_WIDTH ), 
.TRIG14_MATCH_TYPE           (FLA1_TRIG14_MATCH_TYPE ), 
.TRIG14_EXCLUDE           (FLA1_TRIG14_EXCLUDE ), 
.TRIG15_PORT_WIDTH           (FLA1_TRIG15_PORT_WIDTH ), 
.TRIG15_MATCH_UNIT            (FLA1_TRIG15_MATCH_UNIT ), 
.TRIG15_CNT_WIDTH           (FLA1_TRIG15_CNT_WIDTH ), 
.TRIG15_MATCH_TYPE           (FLA1_TRIG15_MATCH_TYPE ), 
.TRIG15_EXCLUDE           (FLA1_TRIG15_EXCLUDE )
) 
u_debug_core_1( 
.drck_in      (drck_o),  
.hub_tdi      (conf_tdi),  
.id_i         (id_o),  
.shift_i      (shift_d), 
.capt_i               (capt_o),  
.conf_sel     (conf_sel[1]),  
.hub_tdo      (hub_tdo[1]),  
.clk          (fla1_clk),  
.resetn_i     (fla1_rstn),  
.trig0_i       (fla1_trig0_i),  
.trig1_i       (fla1_trig1_i),  
.trig2_i       (fla1_trig2_i),  
.trig3_i       (fla1_trig3_i),  
.trig4_i       (fla1_trig4_i),  
.trig5_i       (fla1_trig5_i),  
.trig6_i       (fla1_trig6_i),  
.trig7_i       (fla1_trig7_i),  
.trig8_i       (fla1_trig8_i),  
.trig9_i       (fla1_trig9_i),  
.trig10_i       (fla1_trig10_i),  
.trig11_i       (fla1_trig11_i),  
.trig12_i       (fla1_trig12_i),  
.trig13_i       (fla1_trig13_i),  
.trig14_i       (fla1_trig14_i),  
.trig15_i       (fla1_trig15_i),  
.data_i       (fla1_data_i)  
); 
endmodule 
