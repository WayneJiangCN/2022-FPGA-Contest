module frame_write_read(

   );
endmodule